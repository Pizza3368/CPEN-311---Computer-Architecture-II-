module datapath(input slow_clock, input fast_clock, input resetb,
                input load_pcard1, input load_pcard2, input load_pcard3,
                input load_dcard1, input load_dcard2, input load_dcard3,
                output [3:0] pcard3_out,
                output [3:0] pscore_out, output [3:0] dscore_out,
                output[6:0] HEX5, output[6:0] HEX4, output[6:0] HEX3,
                output[6:0] HEX2, output[6:0] HEX1, output[6:0] HEX0);
						
// The code describing your datapath will go here.  Your datapath 
// will hierarchically instantiate six card7seg blocks, two scorehand
// blocks, and a dealcard block.  The registers may either be instatiated
// or included as sequential always blocks directly in this file.
//
// Follow the block diagram in the Lab 1 handout closely as you write this code.
	// module dealcard(input clock, input resetb, output [3:0] new_card);
	// module card7seg(input [3:0] card, output[6:0] seg7);
	//module scorehand(input [3:0] card1, input [3:0] card2, input [3:0] card3, output [3:0] total);
	reg[3:0] newcard;
	reg[3:0] playercard1;
	reg[3:0] playercard2;
	reg[3:0] playercard3;
	reg[3:0] dealercard1;
	reg[3:0] dealercard2;
	reg[3:0] dealercard3;
	
	// dealcard generates the random card value and stores it in new card.
	dealcard randomCardGenerator (.clock(fast_clock), .resetb(resetb), .new_card(newcard));
	
	// newcard is connected to the 6 registers below:
	// Player registers: Stores playcards in playercard1, playercard2, playercard3.
	reg4 player1_register(.in(newcard), .reset(resetb), .clock(slow_clock), .enabled(load_pcard1), .out(playercard1));
	reg4 player2_register(.in(newcard), .reset(resetb), .clock(slow_clock), .enabled(load_pcard2), .out(playercard2));
	reg4 player3_register(.in(newcard), .reset(resetb), .clock(slow_clock), .enabled(load_pcard3), .out(playercard3));

	// Dealer registers: Stores dealercards in dealercard1, dealercard2, dealercard3.
	reg4 dealer1_register(.in(newcard), .reset(resetb), .clock(slow_clock), .enabled(load_dcard1), .out(dealercard1));
	reg4 dealer2_register(.in(newcard), .reset(resetb), .clock(slow_clock), .enabled(load_dcard2), .out(dealercard2));
	reg4 dealer3_register(.in(newcard), .reset(resetb), .clock(slow_clock), .enabled(load_dcard3), .out(dealercard3));

	// All the outputs of the registers are connected to the card7seg which outputs Hex that are shows the number on the 7 segment LED.
	// player card 1 LED:
	card7seg led_player1(.card(playercard1), .seg7(HEX0));

	// player card2 LED:
	card7seg led_player2(.card(playercard2), .seg7(HEX1));

	// player card3 LED:
	card7seg led_player3(.card(playercard3), .seg7(HEX2));

	// dealer card1 LED:
	card7seg led_dealer1(.card(dealercard1), .seg7(HEX3));

	// dealer card2 LED:
	card7seg led_dealer2(.card(dealercard2), .seg7(HEX4));

	// dealer card3 LED:
	card7seg led_dealer3(.card(dealercard3), .seg7(HEX5));

	// Player card 1,2,3 are used to calculate the current score of player using the scorehand module:
	scorehand player_sch(.card1(playercard1), .card2(playercard2), .card3(playercard3), .total(pscore_out));

	// dealer card 1,2,3 are used to calculate the current score of dealer using the scorehand module:
	scorehand delaer_sch(.card1(dealercard1), .card2(dealercard2), .card3(dealercard3), .total(dscore_out));

	// we need assign whatever the value of player card3 in pcard3_out. 
	assign pcard3_out = playercard3;
	
endmodule

module reg4(input [3:0] in, input reset, input clock, input enabled, output [3:0] out);
	reg[3:0] outvalue;
	// synchronous reset (active-low)
	always @(posedge clock) 
		begin
			if (reset == 0) begin
				outvalue = 4'b0000;
			end
			else begin
				 if (enabled == 1) begin
					outvalue = in;
				end
				// nothing when enabled is 0, keep the old value. 
			end
		end
	assign out =  outvalue;
endmodule