`define startk 4'b0000
`define readi 4'b0001
`define savei 4'b0010
`define modifyj 4'b0011
`define readj 4'b0100
`define savej 4'b0101
`define writei 4'b0110
`define writej 4'b0111
`define incrementi 4'b1000
`define finishk 4'b1001

/* Essentially writing to S. */
// addr, wrdata, wren, rdy
module ksa(input logic clk, input logic rst_n,
           input logic en, output logic rdy,
           input logic [23:0] key,
           output logic [7:0] addr, input logic [7:0] rddata, output logic [7:0] wrdata, output logic wren);

    reg [7:0] i = 8'd0; /* i-th index */
    reg[7:0] j = 8'd0; /* j-th index */

    reg[7:0] valuei = 8'd1; /* value of s[i] */
    reg[7:0] valuej = 8'd1; /* value of s[j] */

    reg finish_flag = 0; /*flag to check if iteration should be done */

    reg[8:0] key_byte = 8'd0;
    reg[3:0] present_state;
    
    always @(posedge clk or negedge rst_n) begin 
        
        if (rst_n == 0) begin
            present_state = `startk; 

            i = 0;
            j = 0;

            rdy = 1;

            wren = 0;
            wrdata = 0;
            addr = 0;
        end

        else begin 
            case (present_state) 

                /* We stay in the start state until enable becomes 1.*/
                `startk: begin 
                    if (en == 1) begin 
                        present_state = `readi;
                    end
                    else begin 
                        present_state = `startk;
                    end
                end

                /* setting s_address to i*/
                `readi: begin 
                    present_state = `savei;
                end

                /* valuei = s[i]*/
                `savei: begin 
                    present_state = `modifyj;
		            valuei = rddata; 
                end

                `modifyj: begin 
                    present_state = `readj;
                    /* key is big endian */
                    case(i % 3)
                        0: key_byte = key[23:16];
                        1: key_byte = key[15:8];
                        2: key_byte = key[7:0];
                        default: key_byte = 8'bx; /*not possible*/
                    endcase
                    j = (j + valuei + key_byte) % 256;
                end

                /* set s address to j
                address = j 8*/
                `readj: begin 
                    present_state = `savej;
		            
                end

                /* valuej = s[j] */
                `savej: begin 
                    present_state = `writei;
                    valuej = rddata;
                end

                // s[i] = s[j]
                // address = j, wren = 1.
                `writei: begin 
                    present_state = `writej;
                end

                // s[j] = s[i]
                `writej: begin 
                    if (finish_flag == 0) begin 
                        present_state = `incrementi;
                    end
                    else begin 
                        present_state = `finishk;
                    end
                end

                // i ++
                `incrementi: begin 
                    present_state = `readi;
                end

                `finishk: begin 
                    if (en == 1) begin 
                        present_state = `readi;
                    end
                    else begin 
                        present_state = `finishk;
                    end
                end

                default: present_state = `startk;
            endcase


            case (present_state) 
                `startk: begin 
                    i = 0;
                    j = 0;
                    rdy = 1;
                    wren = 0;
                    addr = 0;
                    wrdata = 0;
                    finish_flag = 0;
                end

                `readi: begin 
                    wrdata = 0;
                    rdy = 0;
                    addr = i; /* read at address i */
                    wren = 0;
                end

                `savei: begin 
                    rdy = 0;
                    wrdata = 0;
                    addr = 0;
                    wren = 0;
                    
                end

                `modifyj: begin
                    rdy = 0;
                    wren = 0;
                    wrdata = 0;
                    wrdata = 0;
                end

                `readj: begin 
                    rdy = 0;
                    addr = j;
                    wren = 0;
                    wrdata = 0;
                end

                `savej: begin 
                    rdy = 0;
                    addr = 0;
                    wren = 0;
                    wrdata = 0;
                end

                `writei: begin 
                    rdy = 0;
                    addr = i;
                    wren = 1;
                    wrdata = valuej;
                end

                /* address = j, wren = 1, wrdata = valuei*/
                `writej: begin 
                    rdy = 0;
                    addr = j;
                    wren = 1;
                    wrdata = valuei;
                end

                `incrementi: begin
                    rdy = 0; 
                    addr = 0;
                    wren = 0;
                    wrdata = 0;
                    i = i+8'd1; // i++
                    if (i == 8'd255) begin 
                        finish_flag = 1;
                    end
                    else begin 
                        finish_flag = 0;
                    end
                end

                `finishk: begin 
			i = 0;
			j = 0;
            finish_flag = 0;
                    addr = 0;
                    rdy = 1;
                    wren = 0;
                    wrdata = 0;
                end

                /*Technically not possible just in case. */
                default: begin 
                    rdy = 0;
                    wren = 0;
                    wrdata = 0;
                    addr = 0;
                end
            endcase
        end
    end


endmodule: ksa
