module tb_datapath();
		reg slow_clock;
		reg fast_clock;
		reg resetb;
		reg load_pcard1;
		reg load_pcard2;
		reg load_pcard3;
		reg load_dcard1;
		reg load_dcard2;
		reg load_dcard3;
		wire[3:0] pcard3_out;
		wire[3:0] pscore_out;
		wire[3:0] dscore_out;
		wire[6:0] HEX5;
		wire[6:0] HEX4;
		wire[6:0] HEX3;
		wire[6:0] HEX2;
		wire[6:0] HEX1;
		wire[6:0] HEX0;

		datapath db(slow_clock, fast_clock, resetb,
                load_pcard1, load_pcard2, load_pcard3,
                load_dcard1, load_dcard2, load_dcard3,
                pcard3_out,
                pscore_out, dscore_out,
                HEX5, HEX4, HEX3,
                HEX2, HEX1, HEX0); 

		always begin
        		#5 slow_clock = ~slow_clock; 
			#15 fast_clock = ~fast_clock;
    		end
		
		// these are used to check if card value changed or not. 
		reg[3:0] p_card1_val;
		reg[3:0] p_card2_val;
		reg[3:0] p_card3_val;
		reg[3:0] d_card1_val;
		reg[3:0] d_card2_val;
		reg[3:0] d_card3_val;
		initial begin
			slow_clock = 0;
			fast_clock = 0;
			resetb = 0;
			load_pcard1 = 0;
			load_pcard2 = 0;
			load_pcard3 = 0;
			load_dcard1 = 0;
			load_dcard2 = 0;
			load_dcard3 = 0;
			#50 // resetb needs to be 0 in the first rising edge of the fast_clock.
			
			resetb = 1; // keep reset at 1.
			#5

			// test load_pcard1.
			load_pcard1 = 1; // only HEXO should show ACE (1) rest of them should be should show BLANK.
			load_pcard2 = 0;
			load_pcard3 = 0;
			load_dcard1 = 0;
			load_dcard2 = 0;
			load_dcard3 = 0;
			#40
			// on the next rising edge of the clock. playercard1 needs to be equal to the random value generated by dealcard.
			if(db.playercard1 != db.newcard) begin $display("Test 1 failed, player card1 is expected to be: %b, actually it is: %b", db.newcard, db.playercard1); end
			// make sure other cards are 0 at this point.
			else if (db.playercard2 != 4'b0000 || db.playercard3 != 4'b0000 || db.dealercard1 != 4'b0000 || db.dealercard2 != 4'b0000 
				|| db.dealercard3 != 4'b000) begin $display("Test 1 failed, other cards are not 0"); end
			else if (pcard3_out != db.playercard3) begin $display("Test 1 failed because pcard3 was not assigned correct value."); end
			else begin $display("Test 1 passed"); end

			// Now set load_dcard1 = 1.
			load_pcard1 = 0;
			load_pcard2 = 0; 
			load_pcard3 = 0;
			load_dcard1 = 1;
			load_dcard2 = 0;
			load_dcard3 = 0;
			p_card1_val = db.playercard1;
			#40
			// on the next rising edge of the clock. playercard1 value should not change to newvalue but dealercard1 should change to new value.
			if (db.playercard1 != p_card1_val || db.dealercard1 != db.newcard) begin $display("Test 2 Failed dealer card1 did not get new value"); end
			// rest of the card should be 0.
			else if (db.playercard2 != 4'b0000 || db.playercard3 != 4'b0000 || db.dealercard2 != 4'b0000 
				|| db.dealercard3 != 4'b000) begin $display("Test 2 failed, other cards are not 0"); end
			else if (pcard3_out != db.playercard3) begin $display("Test 2 failed because pcard3 was not assigned correct value."); end
			else begin $display("Test 2 passed"); end
			

			// Now set load_pcard2 = 1.
			load_pcard1 = 0;
			load_pcard2 = 1; 
			load_pcard3 = 0;
			load_dcard1 = 0;
			load_dcard2 = 0;
			load_dcard3 = 0;
			d_card1_val = db.dealercard1;
			#40
			// on the next rising edge of the clock, playercard2 should get newcard but playercard1 and dealercard should not change.
			if (db.playercard1 != p_card1_val || db.dealercard1 != d_card1_val || db.playercard2 != db.newcard) begin
			$display("Test 3 failed on first case");
			end
			// check if other registers are 0. 
			else if (db.playercard3 != 4'b0000 || db.dealercard2 != 4'b0000 
				|| db.dealercard3 != 4'b000) begin $display("Test 3 failed, other cards are not 0"); end
			else if (pcard3_out != db.playercard3) begin $display("Test 3 failed because pcard3 was not assigned correct value."); end
			else begin $display("Test 3 passed"); end

			// Now set load_dcard2 = 1. 
			load_pcard1 = 0;
			load_pcard2 = 0; 
			load_pcard3 = 0;
			load_dcard1 = 0;
			load_dcard2 = 1;
			load_dcard3 = 0;
			p_card2_val = db.playercard2;
			#40
			// on the next rising edge of the clock, dealer card2 shoudl get new card but player card1,2 and dealer card1 shoud remain the same.
			if (db.playercard1 != p_card1_val || db.playercard2 != p_card2_val || db.dealercard1 != d_card1_val || db.dealercard2 != db.newcard) begin
			$display("Test 4 failed on first case");
			end
			// check if other registers are 0. 
			else if (db.playercard3 != 4'b0000 
				|| db.dealercard3 != 4'b000) begin $display("Test 4 failed, other cards are not 0"); end
			else if (pcard3_out != db.playercard3) begin $display("Test 5 failed because pcard3 was not assigned correct value."); end
			else begin $display("Test 4 passed"); end

			// now set load_pcard3 = 1.
			load_pcard1 = 0;
			load_pcard2 = 0; 
			load_pcard3 = 1;
			load_dcard1 = 0;
			load_dcard2 = 0;
			load_dcard3 = 0;
			d_card2_val = db.dealercard2;
			#40
			// on next risign edge of the clock, playercard3 will get new value, playercard1, 2 should hold old value
			// dealercard1, 2 should hold the old value.
			if (db.playercard1 != p_card1_val || db.playercard2 != p_card2_val || db.dealercard1 != d_card1_val || db.dealercard2 != d_card2_val
				|| db.playercard3 != db.newcard) begin
			$display("Test 5 failed on first case");
			end
			// check if other registers are 0. 
			else if (db.dealercard3 != 4'b000) begin $display("Test 5 failed, other cards are not 0"); end
			// check if pcard3_out gets the correct value.
			else if (pcard3_out != db.playercard3) begin $display("Test 5 failed because pcard3 was not assigned correct value."); end
			else begin $display("Test 5 passed"); end

			// now set load_dcard3 = 1
			load_pcard1 = 0;
			load_pcard2 = 0; 
			load_pcard3 = 0;
			load_dcard1 = 0;
			load_dcard2 = 0;
			load_dcard3 = 1;
			p_card3_val = db.playercard3;
			#40
			// on next rising edge of the clock, dealer card3 should get new value, playercard 1,2,3 should hold old value and
			// dealer card 1,2 should hold old value. 
			if (db.playercard1 != p_card1_val || db.playercard2 != p_card2_val || db.playercard3 != p_card3_val || db.dealercard1 != d_card1_val 
				|| db.dealercard2 != d_card2_val
				|| db.dealercard3 != db.newcard) begin
			$display("Test 6 failed on first case");
			end
			else if (pcard3_out != db.playercard3) begin $display("Test 5 failed because pcard3 was not assigned correct value."); end
			else begin $display("Test 6 passed"); end
			
			// Now set all of them to 0.
			load_pcard1 = 0;
			load_pcard2 = 0; 
			load_pcard3 = 0;
			load_dcard1 = 0;
			load_dcard2 = 0;
			load_dcard3 = 0;
			d_card3_val = db.dealercard3;
			#40
			// on next risign edge of the clock, all playercard should hold old value. 
			if (db.playercard1 != p_card1_val || db.playercard2 != p_card2_val || db.playercard3 != p_card3_val || db.dealercard1 != d_card1_val 
				|| db.dealercard2 != d_card2_val
				|| db.dealercard3 != d_card3_val) begin
			$display("Test 7 failed on first case");
			end
			else if (pcard3_out != db.playercard3) begin $display("Test 7 failed because pcard3 was not assigned correct value."); end
			else begin $display("Test 7 passed"); end

			// set reset to 0: basically showing a restart of game.
			// this should make all player cards and dealer cards to be 0.
			resetb = 0;
			#40 // wait for next clock cycle.
			if (db.playercard1 != 4'b0000 || db.playercard2 != 4'b0000 || db.playercard3 != 4'b0000 || db.dealercard1 != 4'b0000 
				|| db.dealercard2 != 4'b0000
				|| db.dealercard3 != 4'b0000) begin
			$display("Test 8 failed. One of the playercards or dealer card was not zero.");
			end
			else if (pcard3_out != db.playercard3) begin $display("Test 8 failed because pcard3 was not assigned correct value."); end
			else begin $display("Test 8 passed"); end	
			
			
		end
		

						
endmodule

