`timescale 1 ps / 1 ps
module tb_rtl_task5();

	reg clk;
	reg [3:0] KEY;
	reg [9:0] SW;
	
	wire [6:0] HEX0;
	wire [6:0] HEX1;
	wire [6:0] HEX2;
	wire [6:0] HEX3;
	wire [6:0] HEX4;
	wire [6:0] HEX5;
	wire [9:0] LEDR;

    task5 t5(
        .CLOCK_50(clk),
        .KEY(KEY),
        .SW(SW),
        .HEX0(HEX0), 
        .HEX1(HEX1), 
        .HEX2(HEX2),
        .HEX3(HEX3), 
        .HEX4(HEX4), 
        .HEX5(HEX5),
        .LEDR(LEDR)
    );

    initial forever begin
        clk = 0;
        #5
        clk = 1;
        #5;
    end

    initial 
    
    begin 

        // write test 1 in CT memory
        $readmemh("D:/Cpen311/Lab-3/Lab-3-CPEN311/task4/test3.memh", 
	        t5.ct.altsyncram_component.m_default.altsyncram_inst.mem_data);
        KEY[3] = 0;
        //SW[9:0] = 10'b0000011000;

        #30
        KEY[3] = 1;

        #1000

	    $display("Done");
    end

endmodule: tb_rtl_task5
